interface spi_intf(input clock);

   logic SCK;
   logic SDI;
   logic SDO;
   logic CSN;
   logic SS;

   logic RESETn;
   
endinterface // spi_intf

   
