package apb_test_pkg;

    `include "uvm_macros.svh"

    import uvm_pkg::*;

    import apb_env_pkg::*;


    `include "apb_base_test.svh"

    `include "apb_init_test.svh"
    `include "apb_reset_test.svh"



endpackage //apb_test_pkg
