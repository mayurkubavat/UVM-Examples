interface my_interface;

   bit clock;

   bit sync_1;
   bit sync_2;

endinterface

