package apb_env_pkg;

    `include "uvm_macros.svh"

    import uvm_pkg::*;


    `include "apb_xtn.svh"

    `include "apb_bridge_config.svh"
    `include "apb_slave_config.svh"

    `include "apb_env_config.svh"

    `include "apb_bridge.svh"
    `include "apb_slave.svh"

    `include "apb_subscriber.svh"

    `include "apb_env.svh"

endpackage //apb_env_pkg
