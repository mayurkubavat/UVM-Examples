interface my_interface;

   bit clock;

   // Signals used for debugging HB in testbench
   bit hb_signal;
   bit hb_event;

endinterface

