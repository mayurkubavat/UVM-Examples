package spi_test_pkg;

	`include "uvm_macros.svh"
	import uvm_pkg::*;


	`include "spi_base_test.svh"

endpackage //spi_test_pkg
