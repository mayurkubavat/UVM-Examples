package apb_env_pkg;

    `include "uvm_macros.svh"

    import uvm_pkg::*;


    `include "apb_xtn.svh"
    `include "reset_xtn.svh"

    `include "apb_bridge_config.svh"
    `include "apb_slave_config.svh"

    `include "apb_env_config.svh"
    `include "apb_seqr.svh"
    `include "reset_seqr.svh"

    `include "apb_bridge_seqs.svh"
    `include "apb_bridge_driver.svh"
    `include "apb_bridge_monitor.svh"
    `include "apb_bridge.svh"

    `include "apb_slave_driver.svh"
    `include "apb_slave_monitor.svh"
    `include "apb_slave.svh"

    
    
    `include "reset_seq.svh"
    `include "reset_driver.svh"
    `include "reset_agent.svh"
    `include "apb_subscriber.svh"

    `include "apb_env.svh"

endpackage //apb_env_pkg
