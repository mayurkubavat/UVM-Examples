interface apb_if(input clock);

endinterface //apb_if

