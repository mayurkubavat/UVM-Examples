class baseInterface extends uvm_object;
   `uvm_object_utils(baseInterface)

   function new(string name = "baseInterface");
      super.new(name);
   endfunction

endclass
