/*****************************************************************
 * Filename: test_pkg.sv
 * Class Name: test_pkg
 * Author: Mayur
 * Creation Date: 6 Aug 2015
 * Completion Date: ___ Aug 2015
 * --------------------------------------------------------------
 * **************************************************************/

package test_pkg;

	`include "uvm_macros.svh"
	import uvm_pkg::*;

	`include "ahb_xtn.svh"
	`include "apb_xtn.svh"

	`include "ahb_agent_config.svh"
	`include "apb_agent_config.svh"
	`include "env_config.svh"
	
	`include "ahb_seqs.svh"
	`include "ahb_sequencer.svh"
	`include "ahb_driver.svh"
	`include "ahb_monitor.svh"
	
	`include "apb_driver.svh"
	`include "apb_monitor.svh"

	`include "ahb_agent.svh"
	`include "apb_agent.svh"
	`include "scoreboard.svh"
	`include "vsequencer.svh"

	`include "env.svh"
	`include "vseqs.svh"

	`include "test_base_lib.svh"

endpackage: test_pkg
