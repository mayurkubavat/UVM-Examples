package interfacePackage;

   `include "uvm_macros.svh"
   import uvm_pkg::*;

   `include "baseInterface.svh"

   `include "sumInterface.svh"
   `include "carryInterface.svh"
   `include "inpInterface.svh"

   `include "myTransaction.svh"
   `include "drvSequence.svh"
   `include "myDriver.svh"
   `include "mySequencer.svh"

endpackage
