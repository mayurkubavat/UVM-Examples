class apb_xtn extends uvm_sequence_item;

    `uvm_object_utils(apb_xtn)

    //
    //Methods
    //

    //Constructor
    function new(string name = "apb_xtn");
        super.new(name);
    endfunction //new

endclass //apb_xtn
